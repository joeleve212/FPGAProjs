module cu_top(
  input clk,              // 100MHz clock
  input rst_n,            // reset button (active low)
  output [7:0] led,       // 8 user controllable LEDs
  input usb_rx,           // USB->Serial input
  output usb_tx,           // USB->Serial output
  input [4:0] io_button,
  output [7:0] io_led0,
  output [7:0] io_led1,
  output [7:0] io_led2,
  input [7:0] io_dip0,
  input [7:0] io_dip1,
  input [7:0] io_dip2,
  output [3:0] io_sel,
  output [7:0] io_seg
  );
  
  wire rst;
  
  // The reset conditioner is used to synchronize the reset signal to the FPGA
  // clock. This ensures the entire FPGA comes out of reset at the same time.
  reset_conditioner reset_conditioner(.clk(clk), .in(!rst_n), .out(rst));
  
  assign led = io_button;
  
  assign usb_tx = usb_rx;  // echo the serial data
    
endmodule

module bcd_oneChar(
  input [3:0] binDig,
  output [7:0] segOut
  );
  
  assign segOut = binDig;
  
  
endmodule